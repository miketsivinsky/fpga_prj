//--------------------------------------------------------------------------------------------------
//      project:       led_blink
//	module:        led_blink
//
//	description:   only for test project organisation and build scripts development
//--------------------------------------------------------------------------------------------------

`ifndef LED_BLINK_SVH
`define LED_BLINK_SVH

`include "cfg_params_generated.svh"

`endif // LED_BLINK_SVH

