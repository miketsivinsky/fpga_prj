//--------------------------------------------------------------------------------------------------
//      project:       slon_ip
//	module:        slon_ip
//
//	description:   test and study xilinx ip workflow
//--------------------------------------------------------------------------------------------------

`ifndef SLON_IP_SVH
`define SLON_IP_SVH

`include "cfg_params_generated.svh"

`endif // SLON_IP_SVH

