//--------------------------------------------------------------------------------------------------
//	module:        prescaler_m
//
//	description:   only for test project organisation and build scripts development
//--------------------------------------------------------------------------------------------------

`ifndef PRESCALER_SVH
`define PRESCALER_SVH

`include "cfg_params_generated.svh"

//******************************************************************************
//******************************************************************************
package prescaler_lib;

//------------------------------------------------------------------------------
//    Settings
//

parameter integer COUNTER_WIDTH   = 32;

endpackage : prescaler_lib


`endif // PRESCALER_SVH

