//--------------------------------------------------------------------------------------------------
//      project:       tq1m
//	module:        tq1m
//
//	description:   based at Harry Zhurov tq1 sdc 'slon'
//--------------------------------------------------------------------------------------------------

`ifndef TQ1M_SVH
`define TQ1M_SVH

`include "cfg_params_generated.svh"

`endif // TQ1M_SVH

